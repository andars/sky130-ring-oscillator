* NGSPICE file created from ring-oscillator.ext - technology: sky130A


* Top level circuit ring-oscillator

X0 node_4 node_3 Vdd Vdd sky130_fd_pr__pfet_01v8 w=840000u l=1.01e+06u
X1 node_1 node_5 GND GND sky130_fd_pr__nfet_01v8 w=990000u l=1.01e+06u
X2 node_2 node_1 GND GND sky130_fd_pr__nfet_01v8 w=990000u l=1.01e+06u
X3 node_5 node_4 Vdd Vdd sky130_fd_pr__pfet_01v8 w=840000u l=1.01e+06u
X4 node_3 node_2 Vdd Vdd sky130_fd_pr__pfet_01v8 w=840000u l=1.01e+06u
X5 node_4 node_3 GND GND sky130_fd_pr__nfet_01v8 w=990000u l=1.01e+06u
X6 node_5 node_4 GND GND sky130_fd_pr__nfet_01v8 w=990000u l=1.01e+06u
X7 node_3 node_2 GND GND sky130_fd_pr__nfet_01v8 w=990000u l=1.01e+06u
X8 node_2 node_1 Vdd Vdd sky130_fd_pr__pfet_01v8 w=840000u l=1.01e+06u
X9 node_1 node_5 Vdd Vdd sky130_fd_pr__pfet_01v8 w=840000u l=1.01e+06u
.end

