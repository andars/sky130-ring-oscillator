magic
tech sky130A
timestamp 1610946282
<< nwell >>
rect 271 410 2592 908
<< nmos >>
rect 451 265 552 364
rect 909 264 1010 363
rect 1365 263 1466 362
rect 1826 263 1927 362
rect 2288 263 2389 362
<< pmos >>
rect 451 432 552 516
rect 909 434 1010 518
rect 1365 432 1466 516
rect 1826 433 1927 517
rect 2288 432 2389 516
<< ndiff >>
rect 293 339 451 364
rect 293 295 351 339
rect 406 295 451 339
rect 293 265 451 295
rect 552 353 719 364
rect 552 285 589 353
rect 617 285 719 353
rect 552 265 719 285
rect 749 336 909 363
rect 749 292 803 336
rect 858 292 909 336
rect 749 264 909 292
rect 1010 349 1175 363
rect 1010 281 1044 349
rect 1072 281 1175 349
rect 1010 264 1175 281
rect 1203 324 1365 362
rect 1203 280 1250 324
rect 1305 280 1365 324
rect 1203 263 1365 280
rect 1466 350 1629 362
rect 1466 282 1509 350
rect 1537 282 1629 350
rect 1466 263 1629 282
rect 1664 330 1826 362
rect 1664 286 1711 330
rect 1766 286 1826 330
rect 1664 263 1826 286
rect 1927 350 2091 362
rect 1927 282 1973 350
rect 2001 282 2091 350
rect 1927 270 2091 282
rect 2125 333 2288 362
rect 2125 289 2186 333
rect 2241 289 2288 333
rect 1927 263 2090 270
rect 2125 263 2288 289
rect 2389 330 2551 362
rect 2389 286 2427 330
rect 2482 286 2551 330
rect 2389 263 2551 286
<< pdiff >>
rect 293 498 451 516
rect 293 454 354 498
rect 409 454 451 498
rect 293 432 451 454
rect 552 500 719 516
rect 552 441 588 500
rect 618 441 719 500
rect 552 432 719 441
rect 749 504 909 518
rect 749 460 807 504
rect 862 460 909 504
rect 749 434 909 460
rect 1010 510 1175 518
rect 1010 451 1044 510
rect 1074 451 1175 510
rect 1010 434 1175 451
rect 1202 504 1365 516
rect 1202 460 1247 504
rect 1302 460 1365 504
rect 1202 432 1365 460
rect 1466 505 1628 516
rect 1466 446 1509 505
rect 1539 446 1628 505
rect 1466 432 1628 446
rect 1664 507 1826 517
rect 1664 463 1715 507
rect 1770 463 1826 507
rect 1664 433 1826 463
rect 1927 508 2090 517
rect 1927 449 1973 508
rect 2003 449 2090 508
rect 1927 433 2090 449
rect 2125 510 2288 516
rect 2125 466 2173 510
rect 2228 466 2288 510
rect 2125 432 2288 466
rect 2389 501 2551 516
rect 2389 457 2427 501
rect 2482 457 2551 501
rect 2389 432 2551 457
<< ndiffc >>
rect 351 295 406 339
rect 589 285 617 353
rect 803 292 858 336
rect 1044 281 1072 349
rect 1250 280 1305 324
rect 1509 282 1537 350
rect 1711 286 1766 330
rect 1973 282 2001 350
rect 2186 289 2241 333
rect 2427 286 2482 330
<< pdiffc >>
rect 354 454 409 498
rect 588 441 618 500
rect 807 460 862 504
rect 1044 451 1074 510
rect 1247 460 1302 504
rect 1509 446 1539 505
rect 1715 463 1770 507
rect 1973 449 2003 508
rect 2173 466 2228 510
rect 2427 457 2482 501
<< psubdiff >>
rect 362 77 529 101
rect 362 36 392 77
rect 485 36 529 77
rect 362 12 529 36
rect 881 74 1021 88
rect 881 26 908 74
rect 980 26 1021 74
rect 881 12 1021 26
rect 1349 81 1489 95
rect 1349 33 1393 81
rect 1465 33 1489 81
rect 1349 19 1489 33
rect 1814 84 1954 95
rect 1814 36 1861 84
rect 1933 36 1954 84
rect 1814 19 1954 36
rect 2309 88 2449 105
rect 2309 40 2350 88
rect 2422 40 2449 88
rect 2309 29 2449 40
<< nsubdiff >>
rect 460 792 543 806
rect 460 725 476 792
rect 524 725 543 792
rect 460 715 543 725
rect 918 785 1008 803
rect 918 732 931 785
rect 992 732 1008 785
rect 918 716 1008 732
rect 1370 781 1460 799
rect 1370 728 1386 781
rect 1447 728 1460 781
rect 1370 712 1460 728
rect 1835 782 1925 799
rect 1835 729 1850 782
rect 1911 729 1925 782
rect 1835 712 1925 729
rect 2287 780 2377 799
rect 2287 727 2301 780
rect 2362 727 2377 780
rect 2287 712 2377 727
<< psubdiffcont >>
rect 392 36 485 77
rect 908 26 980 74
rect 1393 33 1465 81
rect 1861 36 1933 84
rect 2350 40 2422 88
<< nsubdiffcont >>
rect 476 725 524 792
rect 931 732 992 785
rect 1386 728 1447 781
rect 1850 729 1911 782
rect 2301 727 2362 780
<< poly >>
rect 451 516 552 568
rect 909 518 1010 568
rect 1365 516 1466 569
rect 1826 517 1927 568
rect 451 407 552 432
rect 451 386 463 407
rect 529 386 552 407
rect 451 364 552 386
rect 909 406 1010 434
rect 2288 516 2389 568
rect 909 385 916 406
rect 982 385 1010 406
rect 909 363 1010 385
rect 1365 406 1466 432
rect 1365 385 1377 406
rect 1443 385 1466 406
rect 451 219 552 265
rect 1365 362 1466 385
rect 1826 406 1927 433
rect 1826 385 1838 406
rect 1904 385 1927 406
rect 1826 362 1927 385
rect 2288 406 2389 432
rect 2288 385 2304 406
rect 2370 385 2389 406
rect 2288 362 2389 385
rect 909 219 1010 264
rect 1365 220 1466 263
rect 1826 219 1927 263
rect 2288 219 2389 263
<< polycont >>
rect 463 386 529 407
rect 916 385 982 406
rect 1377 385 1443 406
rect 1838 385 1904 406
rect 2304 385 2370 406
<< locali >>
rect 295 809 2548 887
rect 295 804 1094 809
rect 295 792 616 804
rect 295 725 476 792
rect 524 725 616 792
rect 295 719 616 725
rect 794 785 1094 804
rect 794 732 931 785
rect 992 732 1094 785
rect 794 724 1094 732
rect 1272 804 2548 809
rect 1272 800 2009 804
rect 1272 781 1563 800
rect 1272 728 1386 781
rect 1447 728 1563 781
rect 1272 724 1563 728
rect 794 719 1563 724
rect 295 715 1563 719
rect 1741 782 2009 800
rect 1741 729 1850 782
rect 1911 729 2009 782
rect 1741 719 2009 729
rect 2187 780 2548 804
rect 2187 727 2301 780
rect 2362 727 2548 780
rect 2187 719 2548 727
rect 1741 715 2548 719
rect 295 615 2548 715
rect 339 498 432 615
rect 339 454 354 498
rect 409 454 432 498
rect 339 441 432 454
rect 572 500 671 515
rect 572 441 588 500
rect 618 441 671 500
rect 782 504 875 615
rect 782 460 807 504
rect 862 460 875 504
rect 782 447 875 460
rect 1029 510 1128 516
rect 1029 451 1044 510
rect 1074 451 1128 510
rect 572 421 671 441
rect 1029 422 1128 451
rect 1228 504 1321 615
rect 1228 460 1247 504
rect 1302 460 1321 504
rect 1228 450 1321 460
rect 1490 505 1589 516
rect 1490 446 1509 505
rect 1539 446 1589 505
rect 1699 507 1792 615
rect 1699 463 1715 507
rect 1770 463 1792 507
rect 1699 450 1792 463
rect 1951 508 2050 516
rect 1490 422 1589 446
rect 1951 449 1973 508
rect 2003 449 2050 508
rect 2152 510 2245 615
rect 2152 466 2173 510
rect 2228 466 2245 510
rect 2152 450 2245 466
rect 2410 501 2506 506
rect 2410 457 2427 501
rect 2482 457 2506 501
rect 1951 422 2050 449
rect 2410 429 2506 457
rect 296 407 551 418
rect 296 385 351 407
rect 404 386 463 407
rect 529 386 551 407
rect 404 385 551 386
rect 296 378 551 385
rect 572 406 1009 421
rect 572 385 916 406
rect 982 385 1009 406
rect 572 380 1009 385
rect 1029 406 1466 422
rect 1029 385 1377 406
rect 1443 385 1466 406
rect 1029 381 1466 385
rect 1490 406 1927 422
rect 1490 385 1838 406
rect 1904 385 1927 406
rect 1490 381 1927 385
rect 1951 406 2388 422
rect 1951 385 2304 406
rect 2370 385 2388 406
rect 1951 381 2388 385
rect 326 339 432 357
rect 326 295 351 339
rect 406 295 432 339
rect 326 190 432 295
rect 572 353 671 380
rect 572 285 589 353
rect 617 285 671 353
rect 572 265 671 285
rect 769 336 875 354
rect 769 292 803 336
rect 858 292 875 336
rect 769 190 875 292
rect 1029 349 1128 381
rect 1029 281 1044 349
rect 1072 281 1128 349
rect 1029 266 1128 281
rect 1228 324 1334 351
rect 1228 280 1250 324
rect 1305 280 1334 324
rect 1228 190 1334 280
rect 1490 350 1589 381
rect 1490 282 1509 350
rect 1537 282 1589 350
rect 1951 350 2050 381
rect 1490 266 1589 282
rect 1690 330 1796 348
rect 1690 286 1711 330
rect 1766 286 1796 330
rect 1690 190 1796 286
rect 1951 282 1973 350
rect 2001 282 2050 350
rect 2410 367 2427 429
rect 2492 367 2506 429
rect 1951 266 2050 282
rect 2158 333 2264 348
rect 2158 289 2186 333
rect 2241 289 2264 333
rect 2158 190 2264 289
rect 2410 330 2506 367
rect 2410 286 2427 330
rect 2482 286 2506 330
rect 2410 274 2506 286
rect 295 100 2548 190
rect 295 91 1080 100
rect 295 77 602 91
rect 295 36 392 77
rect 485 36 602 77
rect 295 -3 602 36
rect 832 74 1080 91
rect 832 26 908 74
rect 980 26 1080 74
rect 832 6 1080 26
rect 1310 96 2548 100
rect 1310 81 1526 96
rect 1310 33 1393 81
rect 1465 33 1526 81
rect 1310 6 1526 33
rect 832 2 1526 6
rect 1756 84 2014 96
rect 1756 36 1861 84
rect 1933 36 2014 84
rect 1756 2 2014 36
rect 2244 88 2548 96
rect 2244 40 2350 88
rect 2422 40 2548 88
rect 2244 2 2548 40
rect 832 -3 2548 2
rect 295 -98 2548 -3
<< viali >>
rect 616 719 794 804
rect 1094 724 1272 809
rect 1563 715 1741 800
rect 2009 719 2187 804
rect 351 385 404 407
rect 2427 367 2492 429
rect 602 -3 832 91
rect 1080 6 1310 100
rect 1526 2 1756 96
rect 2014 2 2244 96
<< metal1 >>
rect 297 809 2539 874
rect 297 804 1094 809
rect 297 719 616 804
rect 794 724 1094 804
rect 1272 804 2539 809
rect 1272 800 2009 804
rect 1272 724 1563 800
rect 794 719 1563 724
rect 297 715 1563 719
rect 1741 719 2009 800
rect 2187 719 2539 804
rect 1741 715 2539 719
rect 297 630 2539 715
rect 286 429 2514 516
rect 286 407 2427 429
rect 286 385 351 407
rect 404 385 2427 407
rect 286 367 2427 385
rect 2492 367 2514 429
rect 286 258 2514 367
rect 302 100 2539 185
rect 302 91 1080 100
rect 302 -3 602 91
rect 832 6 1080 91
rect 1310 96 2539 100
rect 1310 6 1526 96
rect 832 2 1526 6
rect 1756 2 2014 96
rect 2244 2 2539 96
rect 832 -3 2539 2
rect 302 -97 2539 -3
<< labels >>
rlabel locali 382 714 382 714 1 Vdd
rlabel locali 447 30 447 30 1 GND
rlabel locali 617 398 617 398 1 node_1
rlabel locali 1058 398 1058 398 1 node_2
rlabel locali 1526 390 1526 390 1 node_3
rlabel locali 1990 398 1990 398 1 node_4
rlabel viali 2447 394 2447 394 1 node_5
<< end >>
